module linalg